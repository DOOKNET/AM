module TOP(
	input	clk,
	input	rst_n,
	output	signed	[15:0]	AM_mod
);





endmodule