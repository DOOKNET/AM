module demodulate(
	input	clk,
	input	rst_n,
	input	
);

endmodule // 