module demodulate(
	input	clk,
	input	rst_n,
	input	signed	[15:0]	AM_mod
);



endmodule
