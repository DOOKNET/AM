module TOP(
	input	sclk,
	input	
);

endmodule // TOP